module registradores (
    input wire [4:0] readRegister1,
    input wire [4:0] readRegister2,
    input wire [4:0] writeRegister,
    input wire [63:0] writeData,
    input wire regWrite,
    input wire clk,
    output reg [63:0] readData1,
    output reg [63:0] readData2
);
    initial begin
        $dumpfile("registers.vcd");
        $dumpvars(0, registradores);
    end
wire [63:0] register0;
wire [63:0] register1;
wire [63:0] register2;
wire [63:0] register3;
wire [63:0] register4;
wire [63:0] register5;
wire [63:0] register6;
wire [63:0] register7;
wire [63:0] register8;
wire [63:0] register9;
wire [63:0] register10;
wire [63:0] register11;
wire [63:0] register12;
wire [63:0] register13;
wire [63:0] register14;
wire [63:0] register15;
wire [63:0] register16;
wire [63:0] register17;
wire [63:0] register18;
wire [63:0] register19;
wire [63:0] register20;
wire [63:0] register21;
wire [63:0] register22;
wire [63:0] register23;
wire [63:0] register24;
wire [63:0] register25;
wire [63:0] register26;
wire [63:0] register27;
wire [63:0] register28;
wire [63:0] register29;
wire [63:0] register30;
wire [63:0] register31;

reg load0;
reg load1;
reg load2;
reg load3;
reg load4;
reg load5;
reg load6;
reg load7;
reg load8;
reg load9;
reg load10;
reg load11;
reg load12;
reg load13;
reg load14;
reg load15;
reg load16;
reg load17;
reg load18;
reg load19;
reg load20;
reg load21;
reg load22;
reg load23;
reg load24;
reg load25;
reg load26;
reg load27;
reg load28;
reg load29;
reg load30;
reg load31;

reg_parametrizado reg0(.clk(clk), .load(1'b1), .in_data(64'd0), .out_data(register0));
reg_parametrizado reg1(.clk(clk), .load(load1), .in_data(writeData), .out_data(register1));
reg_parametrizado reg2(.clk(clk), .load(load2), .in_data(writeData), .out_data(register2));
reg_parametrizado reg3(.clk(clk), .load(load3), .in_data(writeData), .out_data(register3));
reg_parametrizado reg4(.clk(clk), .load(load4), .in_data(writeData), .out_data(register4));
reg_parametrizado reg5(.clk(clk), .load(load5), .in_data(writeData), .out_data(register5));
reg_parametrizado reg6(.clk(clk), .load(load6), .in_data(writeData), .out_data(register6));
reg_parametrizado reg7(.clk(clk), .load(load7), .in_data(writeData), .out_data(register7));
reg_parametrizado reg8(.clk(clk), .load(load8), .in_data(writeData), .out_data(register8));
reg_parametrizado reg9(.clk(clk), .load(load9), .in_data(writeData), .out_data(register9));
reg_parametrizado reg10(.clk(clk), .load(load10), .in_data(writeData), .out_data(register10));
reg_parametrizado reg11(.clk(clk), .load(load11), .in_data(writeData), .out_data(register11));
reg_parametrizado reg12(.clk(clk), .load(load12), .in_data(writeData), .out_data(register12));
reg_parametrizado reg13(.clk(clk), .load(load13), .in_data(writeData), .out_data(register13));
reg_parametrizado reg14(.clk(clk), .load(load14), .in_data(writeData), .out_data(register14));
reg_parametrizado reg15(.clk(clk), .load(load15), .in_data(writeData), .out_data(register15));
reg_parametrizado reg16(.clk(clk), .load(load16), .in_data(writeData), .out_data(register16));
reg_parametrizado reg17(.clk(clk), .load(load17), .in_data(writeData), .out_data(register17));
reg_parametrizado reg18(.clk(clk), .load(load18), .in_data(writeData), .out_data(register18));
reg_parametrizado reg19(.clk(clk), .load(load19), .in_data(writeData), .out_data(register19));
reg_parametrizado reg20(.clk(clk), .load(load20), .in_data(writeData), .out_data(register20));
reg_parametrizado reg21(.clk(clk), .load(load21), .in_data(writeData), .out_data(register21));
reg_parametrizado reg22(.clk(clk), .load(load22), .in_data(writeData), .out_data(register22));
reg_parametrizado reg23(.clk(clk), .load(load23), .in_data(writeData), .out_data(register23));
reg_parametrizado reg24(.clk(clk), .load(load24), .in_data(writeData), .out_data(register24));
reg_parametrizado reg25(.clk(clk), .load(load25), .in_data(writeData), .out_data(register25));
reg_parametrizado reg26(.clk(clk), .load(load26), .in_data(writeData), .out_data(register26));
reg_parametrizado reg27(.clk(clk), .load(load27), .in_data(writeData), .out_data(register27));
reg_parametrizado reg28(.clk(clk), .load(load28), .in_data(writeData), .out_data(register28));
reg_parametrizado reg29(.clk(clk), .load(load29), .in_data(writeData), .out_data(register29));
reg_parametrizado reg30(.clk(clk), .load(load30), .in_data(writeData), .out_data(register30));
reg_parametrizado reg31(.clk(clk), .load(load31), .in_data(writeData), .out_data(register31));


// como o sinal tem so 1 load, precisa ter o load para o registrador
// especifico somente
always @(writeRegister) begin
    if (regWrite == 1) begin
        case (writeRegister)

            5'b0 : begin 
                load0 <= 1'b1;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1 : begin 
                load0 <= 1'b0;
                load1 <= 1'b1;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h2 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b1;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h3 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b1;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h4 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b1;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h5 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b1;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h6 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b1;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h7 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b1;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h8 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b1;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h9 : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b1;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hA : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b1;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hB : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b1;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hC : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b1;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hD : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b1;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hE : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b1;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'hF : begin 
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b1;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h10: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b1;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h11: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b1;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h12: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b1;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h13: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b1;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h14: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b1;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h15: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b1;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h16: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b1;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h17: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b1;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h18: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b1;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h19: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b1;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1A: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b1;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1B: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b1;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1C: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b1;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1D: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b1;
                load30 <= 1'b0;
                load31 <= 1'b0;
            end
            5'h1E: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b1;
                load31 <= 1'b0;
            end
            5'h1F: begin
                load0 <= 1'b0;
                load1 <= 1'b0;
                load2 <= 1'b0;
                load3 <= 1'b0;
                load4 <= 1'b0;
                load5 <= 1'b0;
                load6 <= 1'b0;
                load7 <= 1'b0;
                load8 <= 1'b0;
                load9 <= 1'b0;
                load10 <= 1'b0;
                load11 <= 1'b0;
                load12 <= 1'b0;
                load13 <= 1'b0;
                load14 <= 1'b0;
                load15 <= 1'b0;
                load16 <= 1'b0;
                load17 <= 1'b0;
                load18 <= 1'b0;
                load19 <= 1'b0;
                load20 <= 1'b0;
                load21 <= 1'b0;
                load22 <= 1'b0;
                load23 <= 1'b0;
                load24 <= 1'b0;
                load25 <= 1'b0;
                load26 <= 1'b0;
                load27 <= 1'b0;
                load28 <= 1'b0;
                load29 <= 1'b0;
                load30 <= 1'b0;
                load31 <= 1'b1;
            end
        endcase
    end else begin
        load0 <= 1'b0;
        load1 <= 1'b0;
        load2 <= 1'b0;
        load3 <= 1'b0;
        load4 <= 1'b0;
        load5 <= 1'b0;
        load6 <= 1'b0;
        load7 <= 1'b0;
        load8 <= 1'b0;
        load9 <= 1'b0;
        load10 <= 1'b0;
        load11 <= 1'b0;
        load12 <= 1'b0;
        load13 <= 1'b0;
        load14 <= 1'b0;
        load15 <= 1'b0;
        load16 <= 1'b0;
        load17 <= 1'b0;
        load18 <= 1'b0;
        load19 <= 1'b0;
        load20 <= 1'b0;
        load21 <= 1'b0;
        load22 <= 1'b0;
        load23 <= 1'b0;
        load24 <= 1'b0;
        load25 <= 1'b0;
        load26 <= 1'b0;
        load27 <= 1'b0;
        load28 <= 1'b0;
        load29 <= 1'b0;
        load30 <= 1'b0;
        load31 <= 1'b0;
    end
    
end

always @(readRegister1, readRegister2) begin
        case (readRegister1)
            5'b0 : readData1 = register0;
            5'h1 : readData1 = register1;
            5'h2 : readData1 = register2;
            5'h3 : readData1 = register3;
            5'h4 : readData1 = register4;
            5'h5 : readData1 = register5;
            5'h6 : readData1 = register6;
            5'h7 : readData1 = register7;
            5'h8 : readData1 = register8;
            5'h9 : readData1 = register9;
            5'hA : readData1 = register10;
            5'hB : readData1 = register11;
            5'hC : readData1 = register12;
            5'hD : readData1 = register13;
            5'hE : readData1 = register14;
            5'hF : readData1 = register15;
            5'h10: readData1 = register16;
            5'h11: readData1 = register17;
            5'h12: readData1 = register18;
            5'h13: readData1 = register19;
            5'h14: readData1 = register20;
            5'h15: readData1 = register21;
            5'h16: readData1 = register22;
            5'h17: readData1 = register23;
            5'h18: readData1 = register24;
            5'h19: readData1 = register25;
            5'h1A: readData1 = register26;
            5'h1B: readData1 = register27;
            5'h1C: readData1 = register28;
            5'h1D: readData1 = register29;
            5'h1E: readData1 = register30;
            5'h1F: readData1 = register31;
            default: readData1 = 32'd0;
        endcase

        case (readRegister2)
            5'h0 : readData2 = register0;
            5'h1 : readData2 = register1;
            5'h2 : readData2 = register2;
            5'h3 : readData2 = register3;
            5'h4 : readData2 = register4;
            5'h5 : readData2 = register5;
            5'h6 : readData2 = register6;
            5'h7 : readData2 = register7;
            5'h8 : readData2 = register8;
            5'h9 : readData2 = register9;
            5'hA : readData2 = register10;
            5'hB : readData2 = register11;
            5'hC : readData2 = register12;
            5'hD : readData2 = register13;
            5'hE : readData2 = register14;
            5'hF : readData2 = register15;
            5'h10: readData2 = register16;
            5'h11: readData2 = register17;
            5'h12: readData2 = register18;
            5'h13: readData2 = register19;
            5'h14: readData2 = register20;
            5'h15: readData2 = register21;
            5'h16: readData2 = register22;
            5'h17: readData2 = register23;
            5'h18: readData2 = register24;
            5'h19: readData2 = register25;
            5'h1A: readData2 = register26;
            5'h1B: readData2 = register27;
            5'h1C: readData2 = register28;
            5'h1D: readData2 = register29;
            5'h1E: readData2 = register30;
            5'h1F: readData2 = register31;
            default: readData2 = 32'd0;
        endcase
    end
endmodule